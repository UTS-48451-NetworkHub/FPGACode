library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tx_fifo is
  port (

  );
end tx_fifo;

architecture arch of tx_fifo is

begin

end architecture arch;
