-- Comment here
