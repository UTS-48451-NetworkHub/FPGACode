COUNT_TEST_8_inst : COUNT_TEST_8 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
