library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity eth_tx_tb_driver is
  port (
    clk    : in  std_logic;
    resetn : in  std_logic;
    enable : in std_logic;
    -- AXI-S interface to eth_tx
    tvalid : out std_logic := '0';
    tready : in  std_logic;
    tlast  : out std_logic := '0';
    tdata  : out std_logic_vector(7 downto 0) := (others => '0')
  );
end entity;

architecture rtl of eth_tx_tb_driver is
  ------------------------------------------------------------------------
  -- Ethernet Packet generated by packet_icmp_gen.py
  ------------------------------------------------------------------------
  constant frame_bytes : natural := 70;
  type rom_t is array (0 to frame_bytes - 1) of std_logic_vector(7 downto 0);
  constant frame_rom : rom_t := (
    x"00",
    x"4C",
    x"BE",
    x"EF",
    x"DE",
    x"AD",
    x"11",
    x"11",
    x"DE",
    x"AD",
    x"BE",
    x"EF",
    x"00",
    x"00",
    x"08",
    x"00",
    x"45",
    x"00",
    x"00",
    x"32",
    x"00",
    x"01",
    x"00",
    x"00",
    x"40",
    x"01",
    x"F7",
    x"4B",
    x"C0",
    x"A8",
    x"01",
    x"2C",
    x"C0",
    x"A8",
    x"01",
    x"02",
    x"08",
    x"00",
    x"E1",
    x"30",
    x"12",
    x"34",
    x"00",
    x"01",
    x"48",
    x"65",
    x"6C",
    x"6C",
    x"6F",
    x"20",
    x"28",
    x"46",
    x"72",
    x"6F",
    x"6D",
    x"20",
    x"46",
    x"50",
    x"47",
    x"41",
    x"29",
    x"21",
    x"21",
    x"21",
    x"00",
    x"FE",
    x"F7",
    x"DA",
    x"26",
    x"1E"
  );

  ------------------------------------------------------------------------
  -- Other Parameters
  ------------------------------------------------------------------------
  -- Constants for timing
  constant CLK_FREQ : natural := 100_000_000; -- 100 MHz
  constant TX_PERIOD : natural := CLK_FREQ;    -- 1 second period
  
  -- Counter for 1-second timing and enable edge detection
  signal timer_count : natural range 0 to TX_PERIOD - 1;
  signal tx_trigger : std_logic;
  signal enable_prev : std_logic;
  signal enable_rising : std_logic;
  
  -- ROM address counter and control signals
  signal rom_addr : natural range 0 to frame_bytes - 1;
  signal tx_active : std_logic;
  signal tx_done : std_logic;
  
  -- Delayed handshake for address increment
  signal handshake_d : std_logic;
    
begin

  -- Enable edge detection and 1-second timer process
  timer_process : process(clk)
  begin
    if rising_edge(clk) then
      if resetn = '0' then
        timer_count <= 0;
        tx_trigger <= '0';
        enable_prev <= '0';
        enable_rising <= '0';
      else
        -- Edge detection for enable
        enable_prev <= enable;
        enable_rising <= enable and not enable_prev;
        
        if enable = '0' then
          timer_count <= 0;
          tx_trigger <= '0';
        else
          if timer_count = TX_PERIOD - 1 then
            timer_count <= 0;
            tx_trigger <= '1';
          else
            timer_count <= timer_count + 1;
            tx_trigger <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -- Transmission control process
  tx_control_process : process(clk)
  begin
    if rising_edge(clk) then
      if resetn = '0' or enable = '0' then
        tx_active <= '0';
        rom_addr <= 0;
        tx_done <= '0';
        handshake_d <= '0';
      else
        -- Delay the handshake by one cycle
        handshake_d <= tx_active and tready;
        
        -- Start transmission on enable rising edge or timer trigger
        if (enable_rising = '1' or tx_trigger = '1') and tx_active = '0' then
          tx_active <= '1';
          rom_addr <= 0;
          tx_done <= '0';
        end if;
        
        -- Advance through ROM one cycle after handshake
        if handshake_d = '1' then
          if rom_addr = frame_bytes - 1 then
            -- Transmission complete
            tx_active <= '0';
            tx_done <= '1';
            rom_addr <= 0;
          else
            -- Next byte
            rom_addr <= rom_addr + 1;
          end if;
        end if;
        
        -- Clear done flag
        if tx_done = '1' then
          tx_done <= '0';
        end if;
      end if;
    end if;
  end process;

  -- Connect outputs
  tvalid <= tx_active;
  tlast <= '1' when (tx_active = '1' and rom_addr = frame_bytes - 1) else '0';
  tdata <= frame_rom(rom_addr) when tx_active = '1' else (others => '0');

end architecture;