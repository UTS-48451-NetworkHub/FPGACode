library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TEN_BASE_RX is
    port (
        DATA_IN : in std_logic
    );
end TEN_BASE_RX;

architecture of TEN_BASE_RX is
    begin

    end
