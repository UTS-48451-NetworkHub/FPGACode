library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tx_fsm is
  port (
    clk : in std_logic -- 100 MHz
  );
end tx_fsm;

architecture arch of tx_fsm is

begin

end architecture arch;