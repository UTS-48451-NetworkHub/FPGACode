library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TEN_BASE_TX is
	port (
		TDp : out std_logic;
		TDn : out std_logic
		);
end TEN_BASE_TX;

architecture of TEN_BASE_TX is begin
begin
	

end